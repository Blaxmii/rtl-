`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.08.2024 13:06:23
// Design Name: 
// Module Name: ha_bhv
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ha_bhv(
    input p,
    input q,
    output sum1,
    output carry1
    );
    
assign sum1=p^q;
assign carry1=p&q;

endmodule
